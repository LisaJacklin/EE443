--Lisa Jacklin
-- EE 443 LAb 4 
-- 2/21/2023

-- Mux 4x4

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX4x4 IS
PORT (x1,x2,x3,x4			:IN STD_LOGIC_VECTOR(3 DOWNTO 0);   --INPUT VALUES FOR THE MUX
		SGN 					:IN STD_LOGIC_VECTOR(1 DOWNTO 0);   -- THIS IS MUX SIGNAL
		Y				  		:BUFFER STD_LOGIC_VECTOR(3 DOWNTO 0)); -- OUTPUT VALUES FOR MUX
END MUX4x4;

ARCHITECTURE MUX4x4_BEHAVIORAL OF MUX4x4 IS 
	
	BEGIN
		-- NOTE THAT THE CONTROL SIGNAL FOR THE MUX IS WITHIN THE PROCESS
			U: PROCESS(SGN) IS
			BEGIN
		
			   IF (SGN = "11") THEN Y <= X4;
			ELSIF (SGN = "10") THEN Y <= X3;
			ELSIF (SGN = "01") THEN Y <= X2;
			ELSIF (SGN = "00") THEN Y <= X1;
			END IF;
			
			END PROCESS;
	
END MUX4x4_BEHAVIORAL;