--Lisa Jacklin
-- EE 443 LAb 4 
-- 2/21/2023

-- REG8x16 using all of the other components

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY REG8x16 IS
	PORT ( D 	:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			 EN, CLK :IN STD_LOGIC;	-- THE SIGNAL AND CLOCK SIGNAL
			 Q 	:OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END REG8x16;

ARCHITECTURE REG8x16_BEHAVIORAL OF REG8x16 IS
	-- 8 TO 16 MULTIPLEXER
	COMPONENT mux8X16 IS
		PORT ( I1, I2, I3, I4, I5, I6, I7, I8	:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
				 SGNL										:IN STD_LOGIC_VECTOR (2 DOWNTO 0);
				 Z											:OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
	END COMPONENT;
	
	--THREE TO EIGHT DECODER FOR READ AND WRITE 
	COMPONENT DCD3x8 IS
		PORT (S	:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
				Q 	:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
	END COMPONENT;
	
	-- 8 BIT REGISTER
	COMPONENT REG8 IS
			PORT (D 			:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			WE, CLK  :IN STD_LOGIC;								--NOTE THAT EN HERE IS THE WE (WRITE ENABLED)
			Q			:OUT STD_LOGIC_VECTOR(7 DOWNTO 0 ));
	END COMPONENT;
	
	BEGIN
	--NEED THREE ADDRESS INPUTS: TWO TO READ AND ONE TO WRITE
	
	
	
	--ONE 16 INPUT DIN[15:0]
	
	--TWO DOUT1[15:0], AND DOUT2[15:0] WHICH ARE THE OUTPUTS FROM THE REGISTER SPECIFIED.
	
	
	
	END REG8x16_BEHAVIORAL;