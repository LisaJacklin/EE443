--Lisa Jacklin
-- EE 443 Lab 6
--DCD5x32.vhd
----------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DCD5x32 IS 
	PORT (DCDIN	:IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			DCDOUT :OUT STD_LOGIC_VECTOR(31 DOWNTO 0));	
END DCD5X32;

ARCHITECTURE DCD5X32_BEHAVIOR OF DCD5X32 IS
	COMPONENT DCD3x8 IS
		PORT (S	:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
				Q 	:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));

	END COMPONENT;
	--TO CONNECT THE VALUES FOR THE MINI DECODERS
	--NOTE THAT THE VECTOR IS LARGE BECAUSE THE OUTPUT IS 5 LARGER THAN THE  INPUT
	SIGNAL INTERN : STD_LOGIC_VECTOR(23 DOWNTO 0);
	
	BEGIN
	--USING SEVERAL PORT MAPS, EACH CHUNK OF THE LARGE ONE WILL BE SEPARATED INTO MANAGEABLE PIECES
	
	D1: DCD3X8 PORT MAP (DCDIN (2 DOWNTO 0), INTERN(7 DOWNTO 0));
	D2: DCD3X8 PORT MAP (DCDIN (4 DOWNTO 2), INTERN(15 DOWNTO 8));
	D3: DCD3X8 PORT MAP (DCDIN (3 DOWNTO 1), INTERN(24 DOWNTO 16));
	
	--NOW, TO SETUP THE ACTUAL OUTPUT FACTORS TO BE OUTPUTS FOR THE 5X32 DECODER
	DCDOUT (31 DOWNTO 24) <= INTERN(24 DOWNTO 16);
	DCDOUT (23 DOWNTO 16) <= INTERN(15 DOWNTO 8);
	DCDOUT (15 DOWNTO 8) <= INTERN(7 DOWNTO 0);
	DCDOUT (7 DOWNTO 0) <= "00000001" WHEN DCDIN = "10000" ELSE "00000000";
	
	
END DCD5X32_BEHAVIOR;