----------------------------------------------------------------------------------
--Lisa Jacklin
-- EE 443 Lab 0
-- 1/24/2022
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



entity DCD3x8 is
--  Port ( );
end DCD3x8;

architecture DCD3x8_behavioral of DCD3x8 is
begin


end DCD3x8_behavioral;
