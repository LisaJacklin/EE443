--Lisa Jacklin
-- EE 443 LAb 6
-- 3/28/2023
--INS_MEM.vhd
---------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY INS_MEM IS
	PORT(
		ADDR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		DOUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END INS_MEM;

ARCHITECTURE INS_MEM_BEHAVIOR OF INS_MEM IS
	TYPE TWODARR IS ARRAY(INTEGER RANGE <>) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	
	COMPONENT DCD5x32 IS 
		PORT(
			DCDIN : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			DCDOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
	END COMPONENT;
		
	COMPONENT DCD3x8 IS
		PORT(
			S : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			Q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	END COMPONENT;
	
	SIGNAL IMEM : TWODARR(0 TO 31);
	SIGNAL RE : STD_LOGIC;
	
BEGIN
	PROCESS(ADDR)
	BEGIN
		IF ADDR(15 DOWNTO 6) = "00000000" THEN
			RE <= '1';
		ELSE
			RE <= '0';
		END IF;
	END PROCESS;
	
	D1: DCD5X32 PORT MAP(ADDR(15 DOWNTO 1), IMEM(31 DOWNTO 0));
	
	PROCESS(RE, IMEM)
	BEGIN
		IF RE = '0' THEN
			DOUT <= (OTHERS => 'Z');
		END IF;
		
		IF RE = '1' THEN
			IMEM(0) <= "0000000000000000";
			IMEM(1) <= "0001000000000000";
			IMEM(2) <= "0010000000000000";
			IMEM(3) <= "0011000000000000";
			IMEM(4) <= "0100000000000000";
			IMEM(5) <= "0101000000000000";
			IMEM(6) <= "0110000000000000";
			IMEM(7) <= "0111000000000000";
			IMEM(8) <= "1000000000000000";
			IMEM(9) <= "1001000000000000";
			IMEM(10) <= "1010000000000000";
			IMEM(11) <= "1011000000000000";
			IMEM(12) <= "1100000000000000";
			IMEM(13) <= "1101000000000000";
			IMEM(14) <= "1110000000000000";
			IMEM(15) <= "1111000000000000";
			IMEM(16) <= "0000000000000000";
			IMEM(17) <= "0000000000000000";
			IMEM(18) <= "0000000000000000";
			IMEM(19) <= "0000000000000000";
		END IF;
		
		DOUT <= IMEM(CONV_INTEGER(ADDR(5 DOWNTO 0)));
		
	END PROCESS;