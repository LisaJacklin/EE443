--Lisa Jacklin
--EE 443 Lab 6
--DCD4x16.vhd
------------------------------------------
