--Lisa Jacklin
-- EE 443 Lab 7
--MUX2x16.vhd
-------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX2X16 IS
	PORT(MUXIN1, MUXIN2	:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		  SIGN	:IN STD_LOGIC;
		  OUTMUX :OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END MUX2X16;

ARCHITECTURE MUX2X16_BEHAVIOR OF MUX2X16 IS
	BEGIN
	
	PROCESS (SIGN, MUXIN1, MUXIN2)
		BEGIN
		
		IF (SIGN = '0') THEN OUTMUX( 15 DOWNTO 0) <= MUXIN1(15 DOWNTO 0);
		ELSIF (SIGN = '1') THEN OUTMUX <= MUXIN2;
		END IF;
		
	END PROCESS;
	
END MUX2X16_BEHAVIOR;