--Lisa Jacklin
-- EE 443 Lab 7
-- Mux2x3
-------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX2X3 IS
	PORT(INPU1, INPU2 :IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			SIGNL2X3		:IN STD_LOGIC;
			OUTPU2X3		:OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END MUX2X3;

ARCHITECTURE MUX2X3_BEHAVIOR OF MUX2X3 IS
	BEGIN
	
	PROCESS(SIGNL2X3, INPU1, INPU2)
		BEGIN
		
		IF (SIGNL2X3 = '0') THEN
			OUTPU2X3 <= INPU1;
		ELSIF (SIGNL2X3 = '1') THEN
			OUTPU2X3 <= INPU2;
		END IF;
		
	END PROCESS;
	
END MUX2X3_BEHAVIOR;