--Lisa Jacklin
-- EE 443 LAb 4 
-- 2/21/2023

-- Mux 8x16 USING MUX4X4 BUILT EARLIER

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX8x16 IS
	PORT ( I1, I2, I3, I4, I5, I6, I7, I8	:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			 SGNL										:IN STD_LOGIC_VECTOR (2 DOWNTO 0);
	       Z											:OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END MUX8x16;

ARCHITECTURE MUX8x16_BEHAVIORAL OF MUX8x16 IS

	COMPONENT MUX4x4 IS
		PORT (x1,x2,x3,x4			:IN STD_LOGIC_VECTOR(3 DOWNTO 0);   --INPUT VALUES FOR THE MUX
			  SGN 					:IN STD_LOGIC_VECTOR(1 DOWNTO 0);   -- THIS IS MUX SIGNAL
			  Y				  		:BUFFER STD_LOGIC_VECTOR(3 DOWNTO 0)); -- OUTPUT VALUES FOR MUX	
	END COMPONENT;
	
	SIGNAL A1, A2: STD_LOGIC_VECTOR (15 DOWNTO 0); --THESE WILL BE THE INTERMEDIATE RESULT FROM THE TWO MUXS G1 AND G2
	
	BEGIN
	--THIS FIRST ONE TAKES THE FIRST FOUR BITS AND GIVE AN OUTPUT
	
		G1: MUX4x4 PORT MAP (I1(3 DOWNTO 0), I2(3 DOWNTO 0), I3(3 DOWNTO 0), I4(3 DOWNTO 0),SGNL(1 DOWNTO 0), A1(3 DOWNTO 0));
		G2: MUX4x4 PORT MAP (I1(7 DOWNTO 4), I2(7 DOWNTO 4), I3(7 DOWNTO 4), I4(7 DOWNTO 4),SGNL(1 DOWNTO 0), A1(7 DOWNTO 4));
		G3: MUX4x4 PORT MAP (I1(11 DOWNTO 8), I2(11 DOWNTO 8), I3(11 DOWNTO 8), I4(11 DOWNTO 8),SGNL(1 DOWNTO 0), A1(11 DOWNTO 8));
		G4: MUX4x4 PORT MAP (I1(15 DOWNTO 12), I2(15 DOWNTO 12), I3(15 DOWNTO 12), I4(15 DOWNTO 12),SGNL(1 DOWNTO 0), A1(15 DOWNTO 12));
	
	-- THIS IS THE BOTTOM SECTION OF THE PORT MAPS
	
		G5: MUX4x4 PORT MAP (I5(3 DOWNTO 0), I6(3 DOWNTO 0), I7(3 DOWNTO 0), I8(3 DOWNTO 0),SGNL(1 DOWNTO 0), A2(3 DOWNTO 0));
		G6: MUX4x4 PORT MAP (I5(7 DOWNTO 4), I6(7 DOWNTO 4), I7(7 DOWNTO 4), I8(7 DOWNTO 4),SGNL(1 DOWNTO 0), A2(7 DOWNTO 4));
		G7: MUX4x4 PORT MAP (I5(11 DOWNTO 8), I6(11 DOWNTO 8), I7(11 DOWNTO 8), I8(11 DOWNTO 8),SGNL(1 DOWNTO 0), A2(11 DOWNTO 8));
		G8: MUX4x4 PORT MAP (I5(15 DOWNTO 12), I6(15 DOWNTO 12), I7(15 DOWNTO 12), I8(15 DOWNTO 12),SGNL(1 DOWNTO 0), A2(15 DOWNTO 12));
		
	-- THIS LAST MUX IS TO GIVE THE RESULTING 16 BIT SOLUTION
	
		G9: MUX4x4 PORT MAP (A1(3 DOWNTO 0), A2(3 DOWNTO 0), "0000","0000" ,SGNL(2 DOWNTO 1), Z(3 DOWNTO 0));
		G10: MUX4x4 PORT MAP (A1(7 DOWNTO 4), A2(7 DOWNTO 4), "0000", "0000",SGNL(2 DOWNTO 1), Z(7 DOWNTO 4));
		G11: MUX4x4 PORT MAP (A1(11 DOWNTO 8), A2(11 DOWNTO 8), "0000", "0000",SGNL(2 DOWNTO 1), Z(11 DOWNTO 8));
		G12: MUX4x4 PORT MAP (A1(15 DOWNTO 12), A2(15 DOWNTO 12), "0000", "0000",SGNL(2 DOWNTO 1), Z(15 DOWNTO 12));

END MUX8x16_BEHAVIORAL;
