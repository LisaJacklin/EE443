--Lisa Jacklin
--EE 443 Lab 6
--SHLONE.vhd
----------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SHLONE IS
	PORT( VALU	:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			OUTP	:OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
	
END SHLONE;

ARCHITECTURE SHLONE_BEHAVIOR OF SHLONE IS 
	BEGIN

--RECOMMENDED TO USE FOR GENERATE...HOW?
--FOR I IN 0 TO 15 GENERATE
	
		OUTP (15 DOWNTO 0) <= VALU (14 DOWNTO 0) & '0';


END SHLONE_BEHAVIOR;