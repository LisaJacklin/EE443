----------------------------------------------------------------------------------
-- Lisa Jacklin
-- EE 443 Lab 0 
-- 1/24/2023
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity module is
--  Port ( );
end module;

architecture module_behavioral of module is
begin


end module_behavioral;
