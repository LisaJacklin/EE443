--Lisa Jacklin
-- EE 443 LAb 0 
-- 1/24/2023

--REG16 using REG8

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY REG16 IS
PORT (D 			:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		EN, CLK  :IN STD_LOGIC;
		Q			:OUT STD_LOGIC_VECTOR(15 DOWNTO 0 ));

END REG16;

ARCHITECTURE REG16_BEHAVIORAL OF REG16 IS

	COMPONENT REG8 IS
		PORT (D 			:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
				EN, CLK  :IN STD_LOGIC;
				Q			:OUT STD_LOGIC_VECTOR(7 DOWNTO 0 ));
	END COMPONENT REG8;
	
	BEGIN
		R1: REG8 PORT MAP (D(7 DOWNTO 0),EN,CLK, Q(7 DOWNTO 0));
		R2: REG8 PORT MAP (D(15 DOWNTO 8),EN,CLK, Q(15 DOWNTO 8));
	
	
END REG16_BEHAVIORAL;