--Lisa Jacklin
-- EE443 Lab 0
-- 1/24/2023

--DCD3x8

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DCD3x8 IS
	PORT (S	:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			Q 	:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));

END DCD3x8;

ARCHITECTURE DCD3x8_BEHAVIORAL OF DCD3x8 IS

	BEGIN 
			Q <= "00000001" WHEN S = "000" ELSE
				  "00000010" WHEN S = "001" ELSE
				  "00000100" WHEN S = "010" ELSE
				  "00001000" WHEN S = "011" ELSE
				  "00010000" WHEN S = "100" ELSE
				  "00100000" WHEN S = "101" ELSE
				  "01000000" WHEN S = "110"ELSE
				  "10000000" WHEN S = "111";

	END DCD3x8_BEHAVIORAL;