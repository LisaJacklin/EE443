LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY INS_MEM IS
    PORT(
        ADDR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        DOUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END ENTITY INS_MEM;

ARCHITECTURE INS_MEM_BEHAVIOR OF INS_MEM IS
    COMPONENT DCD5x32 IS 
        PORT(
            DCDIN : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
            DCDOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
        );
    END COMPONENT;
        
    COMPONENT DCD3x8 IS
        PORT(
            S : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            Q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
        );
    END COMPONENT;
    
    TYPE TDARR IS ARRAY(0 to 31) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	 
    SIGNAL IMEM : TDARR(0 TO 31) := (
        0 => X"0000000000000000",   -- Initialize IMEM with desired values
        1 => X"0000000000000000",
        2 => X"0000000000000000",
        3 => X"0000000000000000",
        4 => X"0000000000000000",
        5 => X"0000000000000000",
        6 => X"0000000000000000",
        7 => X"0000000000000000",
        8 => X"0000000000000000",
        9 => X"0000000000000000",
        10 => X"0000000000000000",
        11 => X"0000000000000000",
        12 => X"0000000000000000",
        13 => X"0000000000000000",
        14 => X"0000000000000000",
        15 => X"0000000000000000",
        16 => X"0000000000000000",
        17 => X"0000000000000000",
        18 => X"0000000000000000",
        19 => X"0000000000000000",
        20 => X"0000000000000000",
        21 => X"0000000000000000",
        22 => X"0000000000000000",
        23 => X"0000000000000000",
        24 => X"0000000000000000",
        25 => X"0000000000000000",
        26 => X"0000000000000000",
        27 => X"0000000000000000",
        28 => X"0000000000000000",
        29 => X"0000000000000000",
        30 => X"0000000000000000",
        31 => X"0000000000000000");

BEGIN
    -- NOTE THAT THE DECODER WILL ONLY DO WORK WHEN ADDR(15 DOWNTO 6) ARE ZERO
    -- NOTE THAT ONLY EVEN MEMORY ADDRESSES ARE USED.
	PROCESS(ADDR) IS
BEGIN
    CASE ADDR(15 DOWNTO 9) IS
        WHEN "000000000" =>
            DOUT <= IMEM(TO_INTEGER(UNSIGNED ADDR(5 DOWNTO 0)));
        WHEN OTHERS =>
            DOUT <= (OTHERS => '0');
    END CASE;
END PROCESS;
END ARCHITECTURE INS_MEM_BEHAVIOR;
