LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY INS_MEM IS
    PORT(
        ADDR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        DOUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END ENTITY INS_MEM;

ARCHITECTURE INS_MEM_BEHAVIOR OF INS_MEM IS
    COMPONENT DCD5x32 IS 
        PORT(
            DCDIN : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
            DCDOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
        );
    END COMPONENT;
        
    COMPONENT DCD3x8 IS
        PORT(
            S : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            Q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
        );
    END COMPONENT;
    
    TYPE TDARR IS ARRAY(0 to 31) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	 
    SIGNAL IMEM : TDARR := (
        0 => "0000001010000010",  -- add R1,R2, R0 
        1 => "0000110100000100",  -- subtract
        2 => "1011011100000110",  --lw
        3 => "1111101110001000",  --sw MAKE CONTROL CHECKS
		  4 => "0100000000000000", --jmp to begining
		  5 =>"0000000000000000",
		 6 =>"0000000000000000",
		7 => "0000000000000000",
		 8 =>"0000000000000000",
		 9 =>"0000000000000000",
		10 => "0000000000000000",
		11 => "0000000000000000",
		12 => "0000000000000000",
		13 => "0000000000000000",
		14 => "0000000000000000",
		15 => "0000000000000000",		
		16 =>"0000000000000000",
		17 =>"0000000000000000",
		18 =>"0000000000000000",
		19 =>"0000000000000000",
		20 =>"0000000000000000",
		21 =>"0000000000000000",
		22 =>"0000000000000000",
		23 =>"0000000000000000",
		24 =>"0000000000000000",
		25 =>"0000000000000000",
		26 =>"0000000000000000",
		27 =>"0000000000000000",
		28 =>"0000000000000000",
		29 =>"0000000000000000",
		30 =>"0000000000000000",
		31 =>"0000000000000000"
       );

BEGIN
    -- NOTE THAT THE DECODER WILL ONLY DO WORK WHEN ADDR(15 DOWNTO 6) ARE ZERO
    -- NOTE THAT ONLY EVEN MEMORY ADDRESSES ARE USED.
	
	--NOTE THAT ERROR CHECKING TO MAKE SURE THERE IS NO ADDRESS OVERFLOW AS WELL
	DOUT <= IMEM((TO_INTEGER(UNSIGNED(ADDR (5 downto 1)))));
	
END ARCHITECTURE INS_MEM_BEHAVIOR;
