--Lisa Jacklin
--EE 443 LAb 9 
-- HexDisplay.vhd
---------------------