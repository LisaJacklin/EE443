--Lisa Jacklin
-- EE 443 LAb 8
--PC.vhdl
-------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PC IS
	PORT (PCNEXT	 		:IN STD_LOGIC_VECTOR(15 DOWNTO 0); --DO YOU NEED THIS INPUT...? THINK YES
			CLK, EN, RST	:IN STD_LOGIC; --CONTROL SIGNALS
			PCOUT 			:OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END PC;

ARCHITECTURE PC_BEHAVIOR OF PC IS
	--SIGNAL PC_INTERN : STD_LOGIC_VECTOR (15 DOWNTO 0);
	CONSTANT INC : INTEGER := 4;
	
	BEGIN
	
	PROCESS(CLK, RST)
		BEGIN
				
			IF RST = '1' 
				THEN pcout <= "0000000000000000";
			ELSIF RISING_EDGE(CLK) AND EN = '1' THEN 
				pcout <= pcnext; -- GIVE AN EDGE OF THE CLOCK TO CHECK
			END IF;
				
		END PROCESS;
			
	--PCOUT <= PC_INTERN;
END PC_BEHAVIOR;