LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY INS_MEM IS
    PORT(
        ADDR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        DOUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END ENTITY INS_MEM;

ARCHITECTURE INS_MEM_BEHAVIOR OF INS_MEM IS
    COMPONENT DCD5x32 IS 
        PORT(
            DCDIN : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
            DCDOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
        );
    END COMPONENT;
        
    COMPONENT DCD3x8 IS
        PORT(
            S : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            Q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
        );
    END COMPONENT;
    
    TYPE TDARR IS ARRAY(0 to 31) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	 
    SIGNAL IMEM : TDARR := (
        0 => "0000001010000010",   -- Initialize IMEM with desired values
        1 => "0000110100000100",
        2 => "0001011100000110",
        3 => "0001101110001000",
        4 => "0010000010001010",
        5 => "0010100110001100",
        6 => "0010111000001110",
        7 => "0011101111010000",
        8 => "0100000010010010",
        9 => "0100110100010100",
        10 => "0101011100010110",
        11 => "0101101110011000",
        12 => "0110000010011010",
        13 => "0110110100011100",
        14 => "0111011100011110",
        15 => "0111101110100000",
        16 => "1000000010100010",
        17 => "1000110100100100",
        18 => "1001011100100110",
        19 => "1001101110101000",
        20 => "1010000010101010",
        21 => "1010110100101100",
        22 => "1011011100101110",
        23 => "1011101110110000",
        24 => "1100000010110010",
        25 => "1100110100110100",
        26 => "1101011100110110",
        27 => "1101101110111000",
        28 => "1110000010111010",
        29 => "1110110100111100",
        30 => "1111011100111110",
        31 => "1111101110000000");

BEGIN
    -- NOTE THAT THE DECODER WILL ONLY DO WORK WHEN ADDR(15 DOWNTO 6) ARE ZERO
    -- NOTE THAT ONLY EVEN MEMORY ADDRESSES ARE USED.
	
	--NOTE THAT ERROR CHECKING TO MAKE SURE THERE IS NO ADDRESS OVERFLOW AS WELL
	DOUT <= IMEM((TO_INTEGER(UNSIGNED(ADDR)) + 4194304)/4);
	
END ARCHITECTURE INS_MEM_BEHAVIOR;
