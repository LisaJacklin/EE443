--Lisa Jacklin
-- EE 443 Lab 5
-- 2/28/2023
--ALU4 CODE
------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ALU4 IS
	PORT (A, B 			:IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			LESS, CIN 	:IN STD_LOGIC;
			SEL			:IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			COUT, OVERFLOW, SET, ZERO	:OUT STD_LOGIC;
			F				:OUT STD_LOGIC_VECTOR (3 DOWNTO 0));
	
	END ALU4;
	
ARCHITECTURE ALU4_BEHAVIOR OF ALU4 IS
--BEFORE DOING ANY OF THE WORK, ALL COMPONENTS CREATED BEFORE THIS MUST BE ADDED AS COMPONENTS
COMPONENT MUX4x4 IS
	PORT (x1,x2,x3,x4			:IN STD_LOGIC_VECTOR(3 DOWNTO 0);   --INPUT VALUES FOR THE MUX
			SGN 					:IN STD_LOGIC_VECTOR(1 DOWNTO 0);   -- THIS IS MUX SIGNAL
			Y				  		:BUFFER STD_LOGIC_VECTOR(3 DOWNTO 0)); -- OUTPUT VALUES FOR MUX
END COMPONENT;

COMPONENT BWOR4 IS
	PORT (O1, O2  :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			U		  :OUT STD_LOGIC_VECTOR(3 DOWNTO 0));	
END COMPONENT;

COMPONENT BWAND4 IS
	PORT ( b1, b2 :in STD_LOGIC_VECTOR (3 DOWNTO 0);
			 F					 :OUT STD_LOGIC_VECTOR (3 DOWNTO 0));
END COMPONENT;

COMPONENT ADD4 IS
	PORT ( X,Y			:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		    CIN			:IN STD_LOGIC;
			 SUM			:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			 COUT			:OUT STD_LOGIC);
END COMPONENT;

COMPONENT PINV4 IS 
	PORT ( INP		:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			 SGNL		:IN STD_LOGIC;
			 INVT		:OUT STD_LOGIC_VECTOR(3 DOWNTO 0));		
END COMPONENT;

--NOTE THAT SIGNALS SHOULD BE USED AT SOME POINT
	SIGNAL MUXOUT,BWOROUT, BWANDOUT, ADDOUT, PINOUTA, PINOUTB,SUB,SLT,OVER : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL CADD, CADD2 :STD_LOGIC;
	
	BEGIN --ARCHITECTURE BEGIN	
		--SO FIRST, MUX SHOULD BE USED TO TAKE AND DO 
		OR4:  	BWOR4 PORT MAP (A, B, BWOROUT);
		AND4: 	BWAND4 PORT MAP (A,B,BWANDOUT);
		AD:   	ADD4 PORT MAP (A, B, CIN, ADDOUT, CADD);
		INVA: 	PINV4 PORT MAP (A, LESS, PINOUTA);
		INVB: 	PINV4 PORT MAP (B, LESS, PINOUTB);
		SUBT: 	ADD4 PORT MAP (A, PINOUTB, CIN, SUB, CADD2);
--	
--	PROCESS (SLT, A, B) IS
--		BEGIN	
--			IF (A <= B) THEN SLT <= A;
--			--ELSIF (A =>B) THEN SLT <= B;
--			--ELSE SLT <= A;
--			END IF;	
--	END PROCESS;	
		
--	PROCESS (A, B, OVER,SEL) IS
--		BEGIN
--			IF (A <= B AND SEL = "100") THEN OVER <= "001";
--			ELSIF (A =>B AND SEL = "010") THEN OVER <= "000";
--			ELSE SLT <= A;
--			END IF;
--	END PROCESS;
--		
	PROCESS(BWOROUT, BWANDOUT, ADDOUT, PINOUTA, PINOUTB,SUB,A,B,SEL) IS
	begin
			IF SEL = "000" THEN F<= BWANDOUT;  --AND
		 ELSIF SEL = "001" THEN F<= BWOROUT; --OR
		 ELSIF SEL =  "010" THEN F<= ADDOUT; --ADD
		 ELSIF SEL =  "100" THEN F<= SUB; --SUB 
	   -- ELSIF SEL =  "110" THEN SET<= SLT; --SET LESS THAN
		 ELSIF SEL =  "111" THEN F<= PINOUTA; --NOT
		 ELSE F <= A;
		 END IF;	  
		 
		 COUT <= CADD OR CADD2;
		 --OVERFLOW <= OVER;
	end process;

			
END ALU4_BEHAVIOR;