--Lisa Jacklin
-- EE 443 Lab 6
--ADD16.vhd
---------------------------------------------
library ieee;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ADD16 IS
	PORT( INA, INB :IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			CAIN		:IN STD_LOGIC;
			ADDOUT	:OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			CAOUT		:OUT STD_LOGIC);
END ADD16;

ARCHITECTURE ADD16_BEHAVIOR OF ADD16 IS
--THE 16 BIT ADDER CONSISTS OF ADD4 PERFORMED IN RIPPLE CARRY
component ADD4 is
	PORT(LHO: IN std_logic_Vector(3 downto 0); -- left hand operand
		 RHO: IN STD_LOGIC_VECTOR(3 downto 0); -- right hand operand
		 C0:  IN STD_LOGIC; -- carry in
		 C4: OUT STD_LOGIC; -- carry out
		 OVERFLOW: OUT STD_LOGIC;             -- if there is overflow (numbers  were to big)
		 R:   OUT STD_LOGIC_VECTOR(3 downto 0)); --output of the adder
	End COMPONENT;

	
	--GOING TO ASSIGN SIGNALS HERE
	SIGNAL COUTS,CO,SUM1,SUM2,overflow   : STD_LOGIC_VECTOR(3 DOWNTO 0);
	
	BEGIN
	--BEGINNING PORTMAPS WHICH TAKE THE FIRST 16 BITS
   A1: ADD4 PORT MAP (INA(3 DOWNTO 0), INB (3 DOWNTO 0), CAIN,overflow(0), COUTS(0), ADDOUT(3 DOWNTO 0) );
   A2: ADD4 PORT MAP (INA(7 DOWNTO 4), INB (7 DOWNTO 4), COUTS(0), overflow(1), COUTS(1), ADDOUT(7 DOWNTO 4) );
	A3: ADD4 PORT MAP (INA (11 DOWNTO 8), INB (11 DOWNTO 8), COUTS(1),overflow(2), COUTS(2), ADDOUT(11 DOWNTO 8));
	A4: ADD4 PORT MAP (INA (15 DOWNTO 12), INB (15 DOWNTO 12), COUTS(2), overflow(3), COUTS(3), ADDOUT (15 DOWNTO 12));
	
	CAOUT <= COUTS(0) AND COUTS(1) AND COUTS(2) AND COUTS(3);
	
END ADD16_BEHAVIOR;