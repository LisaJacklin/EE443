LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY INS_MEM IS
    PORT(
        ADDR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        DOUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END ENTITY INS_MEM;

ARCHITECTURE INS_MEM_BEHAVIOR OF INS_MEM IS
    COMPONENT DCD5x32 IS 
        PORT(
            DCDIN : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
            DCDOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
        );
    END COMPONENT;
        
    COMPONENT DCD3x8 IS
        PORT(
            S : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            Q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
        );
    END COMPONENT;
    
    TYPE TDARR IS ARRAY(0 to 4) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	 
    SIGNAL IMEM : TDARR := (
        0 => "0000001010000010",  -- add R1,R2, R0 
        1 => "0001110100000100",  -- subtract
        2 => "1101011100000110",  --lw
        3 => "1101101110001000",  --sw
		  4 => "0100000000000000" --jmp to begining
       );

BEGIN
    -- NOTE THAT THE DECODER WILL ONLY DO WORK WHEN ADDR(15 DOWNTO 6) ARE ZERO
    -- NOTE THAT ONLY EVEN MEMORY ADDRESSES ARE USED.
	
	--NOTE THAT ERROR CHECKING TO MAKE SURE THERE IS NO ADDRESS OVERFLOW AS WELL
	DOUT <= IMEM((TO_INTEGER(UNSIGNED(ADDR)) + 4194304)/4);
	
END ARCHITECTURE INS_MEM_BEHAVIOR;
