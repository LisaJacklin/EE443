--Lisa Jacklin
--EE 443 Lab 5
-- 2/28/2023
--PINV4
-----------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PINV4 IS 
	PORT ( INP		:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			 SGNL		:IN STD_LOGIC;
			 INVT		:OUT STD_LOGIC_VECTOR(3 DOWNTO 0));	
	
END PINV4;

ARCHITECTURE PINV4_BEHAVIORAL OF PINV4 IS
	BEGIN
	I:
	PROCESS (SGNL) IS
		BEGIN
		--THIS SHOULD BE ABLE TO DISPLAY THE INVERSION IF THE SIGNAL IS A SPECIFIED SENSITIVITY
			IF (SGNL = '1') THEN
				INVT <= NOT INP; -- THIS SHOULD INVERT ALL VALUES IN THE INPUT
			ELSE
				INVT <= INP;
			END IF;
	END PROCESS;
	
	
END PINV4_BEHAVIORAL;