--Lisa Jacklin
--EE 443 Lab 6
--SGNEXT6x16.vhd
------------------------------------------