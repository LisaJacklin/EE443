--Lisa Jacklin
-- EE 443 Lab 5
-- 2/28/2023
--ALU4 CODE
------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ALU4 IS
	PORT (A, B 			:IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			LESS, CIN 	:IN STD_LOGIC;
			SEL			:IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			COUT, OVERFLOW, SET, ZERO	:OUT STD_LOGIC;
			F				:OUT STD_LOGIC_VECTOR (3 DOWNTO 0));
	
	END ALU4;
	
ARCHITECTURE ALU4_BEHAVIOR OF ALU4 IS
--BEFORE DOING ANY OF THE WORK, ALL COMPONENTS CREATED BEFORE THIS MUST BE ADDED AS COMPONENTS
COMPONENT MUX4x4 IS
	PORT (x1,x2,x3,x4			:IN STD_LOGIC_VECTOR(3 DOWNTO 0);   --INPUT VALUES FOR THE MUX
			SGN 					:IN STD_LOGIC_VECTOR(1 DOWNTO 0);   -- THIS IS MUX SIGNAL
			Y				  		:BUFFER STD_LOGIC_VECTOR(3 DOWNTO 0)); -- OUTPUT VALUES FOR MUX
END MUX4x4;

COMPONENT BWOR4 IS
	PORT (O1, O2  :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			U		  :OUT STD_LOGIC_VECTOR(3 DOWNTO 0));	
END BWOR4;

COMPONENT BWAND4 IS
	PORT ( b1, b2 :in STD_LOGIC_VECTOR (3 DOWNTO 0);
			 F					 :OUT STD_LOGIC_VECTOR (3 DOWNTO 0));
END BWAND4;

COMPONENT ADD4 IS
	PORT ( X,Y			:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		    CIN			:IN STD_LOGIC;
			 SUM			:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			 COUT			:OUT STD_LOGIC);
END ADD4;

--NOTE THAT SIGNALS SHOULD BE USED AT SOME POINT

	BEGIN
	
	--NOTE THAT MUX4X4 IS TO SELECT ALU OUTPUT BASED ON THE SEL SIGNALS; 
	--A PROCESS WILL BE USED TO SEND OUT THE RESULT F AND OTHER OUTPUT SIGNALS.
	
	--SINCE (SEL) IS THE SIGNAL FOR OPERATION, THERE SHOULD BE A PROCESS
	PROCESS (SEL) IS
		BEGIN 
		
	END PROCESS;
	
	
	
	
	END ALU4_BEHAVIOR;