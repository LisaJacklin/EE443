--Lisa Jacklin
--EE 443 LAb 6
--INCTWO.vhd
-----------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY INCTWO IS
	PORT (INCIN	:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			INCOUT : OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END INCTWO;

ARCHITECTURE INCTWO_BEHAVIOR OF INCTWO IS
	COMPONENT ADD16 IS --IS THIS ADDITION TRULY NEEDED WHEN THE ADDER CAN ONLY OUTPUT 4 BITS?
		PORT( INA, INB :IN STD_LOGIC_VECTOR(15 DOWNTO 0);
				CAIN		:IN STD_LOGIC;
				ADDOUT	:OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
				CAOUT		:OUT STD_LOGIC);
	END COMPONENT;
	 
	 SIGNAL CAO,CIN :STD_LOGIC;
	 
	BEGIN
	
	A1: ADD16 PORT MAP (INCIN(15 DOWNTO 0), X"0002", CIN,INCOUT(15 DOWNTO 0), CAO);
	
	
END INCTWO_BEHAVIOR;