--Lisa Jacklin
--EE 443 Lab 5
--2/28/2023
--ADD4.vhdl
----------------------------------------------

library ieee;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ADD4 IS
	PORT ( X,Y			:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		    CIN			:IN STD_LOGIC;
			 SUM			:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			 COUT			:OUT STD_LOGIC);
	END ADD4;
	
ARCHITECTURE ADD4_BEHAVIORAL OF ADD4 IS
	
	--DO i NEED TO HAVE SIGNALS?
	SIGNAL C1,C2,C3,c4,S1,S2,S3,S4,N1,N2,N3,N4 :STD_LOGIC;
	
	BEGIN
	
	--THESE ARE THE SETS OF RESULTS THAT WILL CARRY THROUGH THE ADDER
	--S REPRESENTS THE NOR GATES AT THE BEGINNING OF EACH GROUP OF BIT 1 AND 1 OF THE TWO VARS
	S1 <=x(0) NOR Y(0);
	S2 <=x(1) NOR Y(1);
	S3 <=x(2) NOR Y(2);
	S4 <=x(3) NOR Y(3);
	
	--N REPRESENTS THE NAND GATES THAT CONNECT THE BITS AS WELL
	N1 <= X(0) NAND Y(0);
	N2 <= X(1) NAND Y(1);
	N3 <= X(2) NAND Y(2);
	N4 <= X(3) NAND Y(3);
	
	--THESE ARE THE INTERMEDIATE CARRY VALUES THAT WILL BE USED TO DETERMINE FINAL SUMS
	C1 <= ((N1) AND CIN) NOR S2 ; --FOR SUM 2
	
	C2 <= (CIN AND N1 AND N2) NOR (N2 AND (S1 OR (NOT S2))); --THE ADDITION OF SEVERAL NOR GATES MAY BE AN ISSUE...
	
	C3 <= ((CIN AND S2 AND S1 AND S3) AND (N2 AND N1 AND S1)) XOR ((N2 AND N1) AND (NOT N2));
	
	C4 <= C3 AND (S4 AND N3) ;
	
	--THESE WILL BE THE RESULTING SUMS
	SUM(0) <= (CIN) XNOR (NOT S1 AND N1);
	
	SUM(1) <= C1 XNOR ((NOT S1) AND N1);
	
	SUM(2) <= C2 XNOR ((NOT S2) AND N2);
	
	SUM(3) <= C3 XNOR ((NOT S3) AND N3);
	
	COUT <= C4 XNOR S4;
	
	END ADD4_BEHAVIORAL;