LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY INS_MEM IS
    PORT(
        ADDR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        DOUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END ENTITY INS_MEM;

ARCHITECTURE INS_MEM_BEHAVIOR OF INS_MEM IS
    COMPONENT DCD5x32 IS 
        PORT(
            DCDIN : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
            DCDOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
        );
    END COMPONENT;
        
    COMPONENT DCD3x8 IS
        PORT(
            S : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            Q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
        );
    END COMPONENT;
    
    TYPE TDARR IS ARRAY(0 to 31) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	 
    SIGNAL IMEM : TDARR(0 TO 31) := (
        0 => X"0000001010000010",   -- Initialize IMEM with desired values
        1 => X"0000110100000100",
        2 => X"0001011100000110",
        3 => X"0001101110001000",
        4 => X"0010000010001010",
        5 => X"0010100110001100",
        6 => X"0010111000001110",
        7 => X"0011101111010000",
        8 => X"0100000010010010",
        9 => X"0100110100010100",
        10 => X"0101011100010110",
        11 => X"0101101110011000",
        12 => X"0110000010011010",
        13 => X"0110110100011100",
        14 => X"0111011100011110",
        15 => X"0111101110100000",
        16 => X"1000000010100010",
        17 => X"1000110100100100",
        18 => X"1001011100100110",
        19 => X"1001101110101000",
        20 => X"1010000010101010",
        21 => X"1010110100101100",
        22 => X"1011011100101110",
        23 => X"1011101110110000",
        24 => X"1100000010110010",
        25 => X"1100110100110100",
        26 => X"1101011100110110",
        27 => X"1101101110111000",
        28 => X"1110000010111010",
        29 => X"1110110100111100",
        30 => X"1111011100111110",
        31 => X"1111101110000000");

BEGIN
    -- NOTE THAT THE DECODER WILL ONLY DO WORK WHEN ADDR(15 DOWNTO 6) ARE ZERO
    -- NOTE THAT ONLY EVEN MEMORY ADDRESSES ARE USED.
	PROCESS(ADDR) IS
BEGIN
    CASE ADDR(15 DOWNTO 9) IS
        WHEN "000000000" =>
            DOUT <= IMEM(TO_INTEGER(STD_LOGIC_VECTOR ADDR(5 DOWNTO 0)));
        WHEN OTHERS =>
            DOUT <= (OTHERS => '0');
    END CASE;
END PROCESS;
END ARCHITECTURE INS_MEM_BEHAVIOR;
