--Lisa Jacklin
--EE 443 Lab 6
--DCD4x16.vhd
------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DCD4X16 IS
	PORT( IN4 :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			CLK :IN STD_LOGIC;
			OUT16 :OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
	
END DCD4X16;

ARCHITECTURE DCD_BEHAVIOR OF DCD4X16 IS
---------COMPONENTS--------------
	COMPONENT DCD3x8 IS
		PORT (S	:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
				Q 	:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
	END COMPONENT;

	SIGNAL INTERMED1, INTERMED2 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	BEGIN
	--GOING TO NEED PORTMAPS TO PULL FOUR TO A SIXTEEN CONVERSION
	D1: DCD3X8 PORT MAP (IN4 (2 DOWNTO 0), INTERMED1);
	
	D2:DCD3X8 PORT MAP (IN4(3)& IN4(1 DOWNTO 0), INTERMED2);
	
	--CONCATINATING THE TWO 3X8 RESULTS
	OUT16 <= INTERMED1 & INTERMED2;
	
END DCD_BEHAVIOR;