--Lisa Jacklin
--EE 443 Lab 6
--INS_MEM.vhd

--find out the propogation delay and resources required for this file and data_mem too
----------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY INS_MEM IS
	PORT(ADDR	:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		  DOUT	:OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
	
END INS_MEM;

ARCHITECTURE INS_MEM_BEHAVIOR OF INS_MEM IS
	TYPE TWODARR IS ARRAY(INTEGER RANGE<>) OF 
			STD_LOGIC_VECTOR (15 DOWNTO 0);
	
	
-------COMPONENTS--------------------------------
	COMPONENT DCD5x32 IS 
		PORT (DCDIN	:IN STD_LOGIC_VECTOR(4 DOWNTO 0);
				DCDOUT :OUT STD_LOGIC_VECTOR(31 DOWNTO 0));	
	END COMPONENT;
		--INCLUDING 3X8 IN ORDER TO TO USE THE 5X32 DECODER
	COMPONENT DCD3x8 IS
	PORT (S	:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			Q 	:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));

	END COMPONENT;
		
	--NOTE THAT THE COLON IN BETWEEN IMEM AND TWO_ADDR IS IMPORTANT! JUST LIKE WHEN USING STD:LOGIC
	--IMEM is for the output of the DCD5x32
	SIGNAL IMEM 	: TWODARR (0 TO 31);
	SIGNAL RE		:STD_LOGIC;
	
	BEGIN
	--NOTE THAT THE DECODER WILL ONLY DO WORK WHEN ADDR(15 DOWNTO 6) ARE ZERO
	--NOTE THAT ONLY EVEN MEMORY ADDRESSES ARE USED.
	PROCESS (ADDR) IS
		BEGIN
			IF (ADDR(15 DOWNTO 6) <= "000000000") THEN RE <= "1";
		   ELSE RE <= "0";
		   END IF;
		END PROCESS;
	
	D1: DCD5X32 PORT MAP (ADDR (5 DOWNTO 1), IMEM(0 TO 31));

	----ASSIGNING MEMORY-------------------------------------

	PROCESS (RE, IMEM) IS
		BEGIN
		
			--FIRST, IF THE RE IS SET TO ZERO, THIS TELL US THERE IS ACCESS ATTEMPT 
			--TO SOMETHING THAT DOESNT EXIST SO IMPEDANCE IS THE OUTPUT
				IF (RE <= "0") THEN DOUT(15 DOWNTO 0) <= "zzzzzzzzzzzzzzzz"; 
			ELSIF RE <= "1" THEN IMEM(0) <= "0000000000000000";
			ELSIF RE <= "1" THEN IMEM(1) <= "";
			ELSIF RE <= "1" THEN IMEM(2) <= "";
			ELSIF RE <= "1" THEN IMEM(3) <= "1000101110101101";
			ELSIF RE <= "1" THEN IMEM(4) <= "";
			ELSIF RE <= "1" THEN IMEM(5) <= "1000101110101101";
			ELSIF RE <= "1" THEN IMEM(6) <= "";
			ELSIF RE <= "1" THEN IMEM(7) <= "";
			ELSIF RE <= "1" THEN IMEM(8) <= "";
			ELSIF RE <= "1" THEN IMEM(9) <= "";
			
			ELSIF RE <= "1" THEN IMEM(10) <= "";
			ELSIF RE <= "1" THEN IMEM(11) <= "";
			ELSIF RE <= "1" THEN IMEM(12) <= "";
			ELSIF RE <= "1" THEN IMEM(13) <= "";
			ELSIF RE <= "1" THEN IMEM(14) <= "";
			ELSIF RE <= "1" THEN IMEM(15) <= "";
			ELSIF RE <= "1" THEN IMEM(16) <= "";
			ELSIF RE <= "1" THEN IMEM(17) <= "";
			ELSIF RE <= "1" THEN IMEM(18) <= "";
			ELSIF RE <= "1" THEN IMEM(19) <= "";
			
			ELSIF RE <= "1" THEN IMEM(20) <= "";
			ELSIF RE <= "1" THEN IMEM(21) <= "";
			ELSIF RE <= "1" THEN IMEM(22) <= "";
			ELSIF RE <= "1" THEN IMEM(23) <= "";
			ELSIF RE <= "1" THEN IMEM(24) <= "";
			ELSIF RE <= "1" THEN IMEM(25) <= "";
			ELSIF RE <= "1" THEN IMEM(26) <= "";
			ELSIF RE <= "1" THEN IMEM(27) <= "";
			ELSIF RE <= "1" THEN IMEM(28) <= "";
			ELSIF RE <= "1" THEN IMEM(29) <= "";
			
			ELSIF RE <= "1" THEN IMEM(30) <= "";
			ELSIF RE <= "1" THEN IMEM(31) <= "";
			
			END IF;
		
		END PROCESS;
			
	
END INS_MEM_BEHAVIOR;