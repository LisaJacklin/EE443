﻿----------------------------------------------------------------------------------
--Lisa Jacklin
-- EE 443 Lab 0
-- 1/24/2022

----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity top is
--  Port ( );
end top;

architecture top_behavioral of top is
begin


end top_behavioral;
